
    `include "apb_base_sequence.sv"
    `include "apb_rd_sequence.sv"
    `include "apb_wr_sequence.sv"
    `include "apb_err_wr_sequence.sv"
    `include "apb_err_rd_sequence.sv"
